    �l  (  0D                o B��� OQ�.�X�/H J�f�"o ��mY�/H #�  dN�  BP�/ N�  �F0< N@NV��//B����    o  � n  h  -f  �X� S� | n  І @Jg  � n  І @H�H��   SgNnj�   Bg0�   Kg,�   Pg,Hy  �BHy  μN�  �LP�Hx��N�  �FX�R�`�R�  �X`�R�  �L`�R�  ��`�R�  �\`�R�  �<`�R���`��   dg��   lg��   sg�`��    o`Hy  �a n /( N�  ��P�#�  �xf* n /( Hy  �cHy  μN�  �L�� Hx N�  �FX�J�  ܈g/9  �xN�  �6X�`
#�  Π  �x�    oR n #�   �|Hy  �v/9  �|N�  ��P�#�  �hf4/9  �|Hy  �xHy  μN�  �L�� Hx N�  �FX�`
#�  ή  �hB�  �(B�  �hN�  �a  �, N�  6F~ #�  ܀N�  : N�  jLN�  jNN�   �J�  �\gHy  ��N�  �X�N�  " N�  .�R�J�  ܀f�J�  �\gHy  ��N�  �X�N�  &�J�  �\gHy  ��N�  �X�N�  '�J�  ܀f�N�  ,:J�f�N�  Sa �/9  �hN�  ��X���  �ho#�  �hJ�f �4/9  �hN�  ��X�J���ga 	�Hx  N�  �FX�,.N^NuNV��H�0�`��(|  �@a �. ���   �-@���   � �   g &n ��   g �   g N�  .$*@�n�� B� /9  �la �X�+@ +y  �P B- B� +L )M y  � (MB� 
�   f Jp` ^N�  .$*@9 .  �Hf$9 L  �IfHy  �Ja BX�+@ � B� `�� B� Hy  �H` �zN�  .$*@� %B-  y  �l .fB( L f: T�/ a �X�+@ ` y  �l -gR�  �l y  �lJf� y  �lJf �B�  - �`�N�  .$*@�n��  y  �l .f( L f T�/ a �X�+@ ` �H y  �l pf ��( c f ��( @ f ��B�  - @ � ` � �   g ���   %g ��   +g �v` �f�   2fB` ���   $f �p L�0�`��N^NuNV��H�8�`��B�  �PB�  �&y  �x(|  �H*L| S�m + R�  @p `
/N�  ��X�. �����g  ��   :fJ�fBp`  ��   
fp��g�B |f<-   f4- l fHm N�  ��X�#�  �P` ��- e f#�     �` �jB |fHy  ��/N�  ��P�J�fp2`N�  |`�   	fR��` �<Bp$L�8�`��N^NuNV��H� �`��*n ~ `�   9n$r
 N�  �bІ�   0. H�H�, �   0l�S�Jg
 -gp ` L� �`��N^NuNV��H�8�`��&y  �B��    g �J�  �\g4+ H�H�/ /+ /+ + H�H�/ H�H�/ Hy  ��N�  ��� H�H��    g ��   g  ��   g N�   $g 2+ H�H�. �   dg�   eg�   ffB+ H�H�+ H�H�၀�, �"<   �N�  �t��  �l(@*T��    g � - ��f LJ�  �\g/ Hy  �N�  �P� g g +f � y  �hS�m ^ y  �hR�  ( S� @� 	p ` R/+ Hy  ��/9  �hN�  �L�� J�  �<g J� g/+ Hy  ��/9  �hN�  �L��  y  �hS�m � y  �hR�  ( S� @� 
p -k ��'y  �( 
#�  �(&n��` �L/9  �h/+ N�  �PP� y  �hS�m y  �hR�  ( S� @� :p `/9  �hHx :N�  ��P�J�  �<g J� g/+ Hy  �/9  �hN�  �L��  y  �hS�m y  �hR�  ( S� @� 
p `/9  �hHx 
N�  ��P�/+ N�  ��X�` �,/9  �hHx 	N�  ��P� y  �hS�m y  �hR�  ( S� @� jp `/9  �hHx jN�  ��P�/9  �h R�/ `@ y  �hS�m y  �hR�  ( S� @� 	p `/9  �hHx 	N�  ��P�/9  �h/N�  �PP��   ff  � y  �hS�m y  �hR�  ( S� @� lp `/9  �hHx lN�  ��P� %f  �/+ /+ Hy  �!/9  �hN�  �L�� J�  �<g J� g/+ Hy  �)/9  �hN�  �L��  y  �hS�m ��` ���   df2 y  �hS�m y  �hR�  ( S� @� b` �`/9  �hHx b` �b�   ef �` y  �hS�m y  �hR�  ( S� @� w` �$/9  �hHx w` �&X���  �He ��(|  �l` ��J� g  � y  �hS�m y  �hR�  ( S� @� 	p `/9  �hHx 	N�  ��P�/9  �h/+ N�  �PP�J�  �<g J� g/+ Hy  �4/9  �hN�  �L��  y  �hS�m ��` �n g g +fd/+ Hy  �?/9  �hN�  �L�� J�  �<g J� g/+ Hy  �E/9  �hN�  �L��  y  �hS�l �\/9  �hHx 
N�  ��P�` �` y  �hS�m�` �8J� gF/9  �h/+ N�  �PP�J�  �<g J� g/+ Hy  �P/9  �hN�  �L�� /+ N�  ��X� y  �hS�m�` ��L�8�`��N^NuNV��H�0�`��*n /N�  ��X�. J�fp `FHx  R�/ N�  �vP�(@��    fHy  �[Hy  μN�  �LP�Hx��aX�//N�  ��P� L�0�`��N^NuNV  J�  �|g/9  �|N�  �X�/. N�  �FX�N^NuNV��/*|  ήJ�  �hg/9  �hHy  �{/N�  �L�� J�  �tg/9  �tHy  ��/N�  �L�� J�  �dg/9  �dHy  ��/N�  �L�� J�  �Tg/9  �THy  ��/N�  �L�� J�  �`g/9  �`Hy  ��/N�  �L�� J�  ��g/9  ��Hy  ��/N�  �L�� J�  ܐg/9  ܐHy  ��/N�  �L�� J�  ܄g/9  ܄Hy  ��/N�  �L�� J�  �8g/9  �8Hy  �/N�  �L�� J�  �g/9  �Hy  �$/N�  �L�� J�  �`g/9  �`Hy  �=/N�  �L�� J�  �pg/9  �pHy  �P/N�  �L�� J�  ܌g/9  ܌Hy  �d/N�  �L�� J�  �Hg/9  �HHy  /N�  �L�� J�  �g/9  �Hy  /N�  �L�� *_N^NuNV��H�8�`��*|  �T`HH�H��+ H�H�Ё�  �"<   �N�  �t��  �d(@`��  �he(|  �dJ�f�Y�(�P�&U��    f�*|  �T`4 �"<   �N�  �t��  �l(@`��  �He(|  �lJ�f�Y�(�P�.- f�L�8�`��N^NuNV��H�< `��&|  ºB+ k  � (|  �H`R� 	g�  g�`  g 	g�Jf�B`R� 	g�  g�#�  �l9  ºH�H��9  »H�H�Ё�  �"<   �N�  �t��  �d$@`j&U(|  º�f
Jf� - `hS�Jf<J, f6 lf - �  f `J bf - �  d `8 wf - �  e `&X���  �he$|  �d*R��    f�#�  �H  �lp L�< `��N^NuNV��H�8 `��&|  ��`B���  ��e�*y  �B`* f "<    - N�  �t��  �� @ �B� *m ��    f�*y  �B`  � g g %g +f  �B� 
"<    - N�  �t��  �� @(P��    g
 - �� g$(y  �B` f
 - �� g(l ��    f��    g./N�  -�X� @-h �� .����g @+h  (n��+L 
R� *m ��    f �N*y  �B`.(m  f"J� f��    gJg %g
/N�  -�X�*L��    f�L�8 `��N^NuNV��H�8 `��B�  ܀*y  �B��    g � g g %fVJ� 
gP/- 
N�  -�X�(@ f<J� g6 - �� g,R�  �t+l  /- 
N�  -�X� l 
R� +l 
 
R�  ܀ fp&m  ff(m 
(l  g���fT/- 
N�  -�X�+k 
 
+k   k !M +k  - H�H��  ¬ @P 'y  �( 
#�  �(R�  ܀R�  �H gv gp`  � m  gh gb g\ $gVJgR !gL "gFR�  ܀R�  �dJ� 
g/( 
N�  -�X�&m  K+h   m !M 'y  �( 
#�  �(J� f�(m ��    gJ fD - 
��fT m !m   m !m  +y  �( 
#�  �(*m /N�  -�X�R�  ܀R�  �T/a&X�/a &X�*@*m ` �*(l `�L�8 `��N^NuNV��H�8 `��*n (m 
��    gd*m ��    g g�(l ��    g g�//N�  ->P�J�g0��g,/a4X�&@� B- +K 
+k  B� R�  ��R�  ܀`�L�8 `��N^NuNV��//(n  g`
(HR�  `T l  g�N�  .$*@� +y  ¶ R�  ¶B� 
B� +|    B� B- +l  +L  l !M )M  (_*_N^NuNV��H�8 `��*n  f (m 
��    fx`  � g| m  f  �(l &L-|   ��&k ��    g  ʷ�g  �S���g  � f� m  + �� f�*m ��    f  � . ` R(l ��    g  � g� f ��(l &m 
`b g fR��gZR�  ܐR�  ܀ m !L  m !K  l !k   k !l  )m  'm  /- 
N�  -�X� `  �&k ��    f� `  ���f �P*n /a �TX�-@��+ H�H��  ¬ @P /+ 
N�  -�X� l !M  k !M  m !L  m !K -m ��+l  )n�� -m ��+k  'n�� /- a ��X�(@'l  'L 
/.��N�  -�X� n��J� nS�  �`R�  �`R�  ܀ L�8 `��N^NuNV��H�8 `��*y  �B`H f>(m 
��    g2�    o(&m ` f + 
��f//a&P�&k ��    f�*m ��    f�L�8 `��N^NuNV��H�< `��*n (n `T/a �X�&@ l !l   l !l  $L(l %y  �( 
#�  �(/, 
N�  -�X�)k  )K 
R�  ܀R�  ܌*m ��    g g�(l //N�  ->P�J�f�L�< `��N^NuNV��H�0�`��*y  �B��    g J�  �\g^~ `D"<   ( N�  �b�  �T @Jg("<   ( N�  �b�  �T/ /Hy  ��N�  ��� R��   m�Hy  ��N�  �X�H�H�S��   -b ��@0; N� ������������B���������������������������������` :Hy  ٬N�  3�X���fX m  gN!m   m !m  +y  �( 
#�  �(R�  �8`  �- e g  �/N�  1�X�Hy  لN�  1�X�. l�Hx Hx  /N�  5 �� Hy  لN�  3�X�. Hy  ٬N�  3�X�, Hy  ٬a 4X�J�mDJ�m"<   ( N�  �b�  �T/ /a ``X/9  ��Hy  ٬N�  9�P�J�fBHy  ٬/`�J�m /9  ��Hy  لN�  9�P�J�fHy  ل`�Hy  ٬Hy  لN�  9HP�Hy  لN�  4�X�*m ` ��- d f ��/N�  1�X�- f fHx Hx  /N�  5 �� Hy  لN�  4�X�Hy  ٬a TX�B9  �,`�/a �X�Hy  لa 8X� f�Hy  لN�  3�X�. mHy  ��/a d`Hy  لHy  ��N�  9HP�`�/a vX�- f fHx  Hx  /N�  5 �� Hy  لN�  4�X�J9  لg �Hy  �,Hy  لN�  9�P�J�g � m !m   m !m  (M*m )y  �( 
#�  �(R�  �R�  ܀` ��/N�  1�X�Hy  ٬N�  4�` � /N�  1�X�Hy  لN�  4�X�Hy  ٬N�  4�X�- f f ��Hy  ٬N�  3�X�J�l<9 #  لf ��Hy  لN�  1�X������f ��Hy  ٬N�  4.X������f ��Hx Hx /N�  5 �� ` �l/N�  6�X�a p` �L�0�`��N^NuNV��H�0�`��~ B���*y  �B`
R�+G *m ��    f�*y  �B`  �(m  f  � f  �J� 
g  ~J� 
gv l 
 , �� / a  �X�-@�� m 
 - �� / ajX�����oF - 
�� 
g<- H�H��  ¬ @P  , 
. )m 
 
+G 
., )m  +G R�  ܄R���*L��    f �^ .��L�0�`��N^NuNV  J� l . D�` . N^NuNV��H�8 `��&n  n �fR+ ( �fFJo m<*k  n (h ��    f ��    g`��    g�fJf�p`
��    f�p L�8 `��N^NuNV��/*n  f.S� n(R�  �` m !m   m !m  +y  �( 
#�  �(*_N^NuNV��/*n `
 f*m ��    f� *_N^NuNV��/*y  �(��    g
#� 
  �(`:Hx  Hx N�  �vP�*@��    f Hy  ��Hy  μN�  �LP�Hx��N�  �X�B- B� B- B� B� 
 *_N^NuNV  B9  ���  ��  פ�  פ  �|�  �|  �TB9  �l�  �l  �D�  �D  ��  �  ��B9  ��  �  ���  ��  ؼ�  ؼ  ؔB9  �\�  �\  �4B9  ��B9  �,N^NuNV��//*n /N�  4�X�J�f&"<   ( . N�  �b�  �T(@�g ,f�S�B(_*_N^NuNV��//~ `J"<   ( N�  �b�  �T*@ af,H�H�". �   (��f"<   ( N�  �b�  �T @BR��   m�.*_N^NuNV��//*n /N�  4�X�/N�  3�X�. m"<   ( N�  �b�  �T @B�   m"/a �RX�`"<   ( N�  �b�  �T @B/N�  1�X�. l� af   0m  � 5n  � @f  �9 #  �TgB9  �T9 #  �|gB9  �|9 #  פgB9  פ9 #  ��gB9  ��9 #  ��gB9  ��9 #  �gB9  �9 #  �DgB9  �D9 #  �lgB9  �l9 #  ؔgB9  ؔ9 #  ؼgB9  ؼ9 #  ��gB9  ��9 #  �gB9  �9 #  �4gB9  �49 #  �\gB9  �\B9  ��.*_N^NuNV��// n *h (|  ل�f�B9  ٬(_*_N^NuNV��H�8 `��&n *k (|  ل` ,g�Jf�B(|  ٬B ,g`R�  g� 	g��f�L�8 `��N^NuNV��/*n Jg �9  �T�f/Hy  �Ta �P�J�gp ` �9  �|�f/Hy  �|a nP�J�gp` �9  פ�f/Hy  פa LP�J�gp` r9  �̰f/Hy  ��a *P�J�gp` P9  ���f/Hy  ��a P�J�gp` .9  ��f/Hy  �a �P�J�gp` 9  �D�f/Hy  �Da �P�J�gp`  �9  �l�f/Hy  �la �P�J�gp`  �9  ؔ�f/Hy  ؔa �P�J�gp`  �9  ؼ�f/Hy  ؼa ^P�J�gp	`  �9  ��f/Hy  ��a <P�J�gp
`b9  ��f/Hy  �a P�J�gp`B9  �4�f/Hy  �4a �P�J�gp`"9  �\�f/Hy  �\a �P�J�gp`p�*_N^NuNV��/*n  df&- 0 m- 7 nJ- f- H�H��   0`. af&- 0 m- 5 nJ- f- H�H��   (`p�*_N^NuNV��/*n  af&- 0 m- 7 nJ- f- H�H��   0` sf- p f
J- fp`p�*_N^NuNV��H�0�`��*n (MJgXJf�, +��g, -��fD af: 0m4 5n.H�H��   (. "<   (N�  �b�  �T @B/N�  /pX�p`p L�0�`��N^NuNV��H�0�`��J� gHy  ٬a ��X�-@��`-|������Hy  لa ��X�. J�lJ���m  �(|  ل*|  ��f�J9  ٬g*|  �<� ,(|  ٬�f�`B9  �<J�mD�   oJ� g  �� a  � �   (`� d  � �   0�  �B9  �R�  �J���mH�   ��oJ� gb� a  �= .���   (`� d  �= .���   0�  �>B9  �?R�  �Hy  �<Hy  �N�  ��P�Hy  �N�  6X� n !@ L�0�`��N^NuNV��//J�  �Bg  �~�*y  �B`l  g !g "fVH�H���gJ� g> m   g !g "f( m !m   m !m  +y  �( 
#�  �(*m `H�H�. *m ��    f�.*_N^NuNV��H�< `��*n (m 
��    g  �/N�  -�X�(@ f/N�  1XX�Hy  �dHx N�  /(P�` f  �/a �HX� l  fn l  g f^Hx adX�&@Hx aZX�$@(l /
/, H�H�/ a  ��� J�g,R�  �pR�  ܀/- 
N�  -�X�+l 
 
+l   m 
R� L�< `��N^NuNV��//"<   ( . N�  �b�  �T*@ #g</a ��X�. m"<   ( N�  �b�  �T`Hy  ��/a zP�J�g <  �` .*_N^NuNV��H�0�`��*n (n  #f  � #f  �~ `  9n r
 N�  �b. H�H��   0ހ 0l�,~ `  9n r
 N�  �b. H�H��   0ހ 0l� +fR� +fR��f  ~Jf� . �   	bl�@0; N�    $ * 0 6 < F P Z`L��fHp`F��f�`>��o�`8��l�`2��m�`,��n�`& "��d`� "��c`� "��b
`� "��d�p L�0�`��N^NuNV��H�8 `��*n (n  #f/aNX�J�g&|  ���f�&|  ��f�L�8 `��N^NuNV��//*n (n �gp `Jf�p(_*_N^NuNV��/*n  *g (g -f- ( fp `Jf�S�S� +g� )fS� 5f�p*_N^NuNV  a 	�N�  t�a N�  t�a �a \aa (a �N^NuNV��H�<�`��*y  �B��    f �` �&l ��    g � f �- f f � f z, f f p f h+ f f ^$k ��    g P f H/N�  1�X�Hy  لN�  3�X�. �   m $�   n Hy  ٬N�  3�X�J�f /N�  1�X�9 #  لf  �Hy  ٬N�  3�X�J�f  �/N�  1�X�Hy  لN�  3�X�J�f  �Hy  ٬N�  4.X�J�f  �/
N�  1�X�9 a  لf  �9 0  مf  �9 @  نf|Hy  ٬N�  3�X�J�fj/N�  1�X�Hy  لHy  �hHn��N�  �Z�� Hn��/a *P�/N�  1�X�Hy  لHy  �nHn��N�  �Z�� Hn��/a �P�/N�  jX�*L(m ��    f �R*y  �B` 4&l ��    g 4 f - f f  f 
, f f   f  �+ f f  �J+ g  �/N�  1�X�Hy  لN�  4.X�. m  ��   n  �Hy  ٬N�  3�X�J�f  �/N�  1�X�9 #  لf  �Hy  ٬N�  3�X�J�f  �/N�  1�X�Hy  لN�  3�X�J�fbHy  ٬N�  4.X���fP/N�  1�X�/Hy  لHy  �tHn��N�  �Z�� Hn��/a �P�//a �P�/N�  jX�/N�  jX�*L(m ��    f ��*y  �B` �&l ��    g � f �- f f � g 
f t, f f j f b+ f f XJ+ g P/N�  1�X�Hy  لN�  3�X�. �   m�   o4Hy  لN�  i|X�J�f"9 _  لg9 .  لf  �9 L  مf  �Hy  ٬N�  3�X�J�f  �/N�  1�X�9 #  لf  �Hy  ٬N�  3�X�J�f  �/N�  1�X�Hy  لN�  3�X�J�f  �Hy  ٬N�  4.X�. m  ��   nx/N�  1�X�/Hy  لHy  �{Hn��N�  �Z�� Hn��/a 2P�/N�  1�X�/Hy  لHy  łHn��N�  �Z�� Hn��/a  P�//a �P�/N�  jX�*L(m ��    f �R*y  �B` V&l ��    g V f >- f f 4 g 
f &, f f  f + f f 
J+ g /N�  1�X�Hy  لN�  4.X�. �����g  �Hy  ٬N�  4.X�J�f  �/N�  1�X�9 #  لf  �Hy  ٬N�  4.X�-@�������g  �/N�  1�X�Hy  لN�  4.X�J�fzHy  ٬N�  4.X�-@�������g`/N�  1�X�����fP����gJ/N�  1�X�/.��Hy  لHy  ŉHn��N�  �Z�� Hn��/a �P�/.��/a �P�/N�  jX�*L(m ��    f ��*y  �B`  f - e f  �J� g  � f  �, f f  �&l ��    g  � f  �+ f f  �/N�  1�X�Hy  ٬N�  3�X�J�f  �/N�  1XX�Hy  لN�  3�X�J�f  �/N�  1�X�Hy  لN�  3�X�J�fjHy  ŐHy  ٬N�  ��P�J�fR/N�  1�X�Hy  لHy  ŕHn��N�  �Z�� Hn��/a zP�/N�  jX�(K� B+ Hy  ś/a XP�*L(m ��    f ��*y  �B` ( f - e f  f , f f &l ��    g  � f  �+ f f  �$k ��    g  �/
N�  ��X�J�g  �/N�  1�X�Hy  ٬N�  3�X�J�f  �/N�  1XX�Hy  لN�  3�X�J�f  �/N�  1�X�Hy  لN�  3�X�J�fjHy  şHy  ٬N�  ��P�J�fR/N�  1�X�Hy  لHy  ŤHn��N�  �Z�� Hn��/a <P�/N�  jX�(K� B+ Hy  Ū/a P�*L(m ��    f ��L�<�`��N^NuNV��/*n *m ��    g  �H�H��   g�   g  �`  �/N�  1�X�Hy  لN�  3�X�J�gHy  لN�  4.X�J�f  �Hy  ٬/. Hy  ŮHn��N�  �Z�� - d fHn��Hy  ŵHy  μN�  �L�� `>Hn��/a LP�`0/N�  1XX�9 a  لf9 0  مf . �   0 m @ *_N^NuNV��H�0�`��*y  �B��    f N` X f g( f g f g f  � f  �- f f  �, f f  �/N�  1�X�Hy  لN�  i|X�J�g  �Hy  ٬N�  3�X�. m  ��   n  �Hy  مN�  h~X�-@��/N�  1�X�Hy  لN�  i|X�J�gfHy  ٬N�  3�X���fTHy  مN�  h~X�Ѯ���   ��n8/N�  jX�Hy  ٬/.��Hy  ��Hn��N�  �Z�� Hn��/a �P�` 0 f g f  f /N�  1�X�Hy  لHn��N�  ��P�Hy  ٬Hn��N�  ��P�/N�  1�X�Hy  ٬Hn��N�  ��P�J�f  �Hn��N�  3�X�. m  �Hy  ٬N�  3�X���f  �- �, f  �Hn��N�  i|X�J�g  �Hy  لN�  i|X�J�glHn��N�  h~X�-@��Hy  مN�  h~X�-@��Hn�� f
 .������` .������/ Hy  ��Hn��N�  �Z�� Hn��/a �P�/N�  jX�(M*L(m ��    f ��L�0�`��N^NuNV��H�8�`��*y  �B��    f �` �- f f  � f  �, f f  �&l ��    g  �J+ g  � f  �J+ g+  g+  g
+  f  �/N�  1�X�Hy  ٬N�  4.X������g|/N�  1�X�Hy  لN�  i|X�J�g`Hy  مN�  h~X�J�fNHy  ٬N�  4.X�. �����g6� /Hy  ��Hn��N�  �Z�� Hn��/a �P�(k `  � g � f  �- f f  � f  �J, g,  g,  g,  frJ, gl/N�  1�X�Hy  لN�  i|X�J�gPHy  مN�  h~X�J�f>Hy  ٬N�  4.X�. �����g&� /Hy  ��Hn��N�  �Z�� Hn��/a 
�P�*L(m ��    f �@L�8�`��N^NuNV��H�< `��*y  �B��    g �(m ��    g Z&l ��    g L f n- d f d f \, e f R f J+ f f @$k ��    g 2 f ** f f  /N�  1�X�Hy  لHn��N�  ��P�Hy  ٬Hn��N�  ��P�/N�  1XX�Hy  لHn��N�  ��P�J�f  �/N�  1XX�Hy  لHn��N�  ��P�J�f  �/
N�  1�X�Hy  ٬Hn��N�  ��P�J�f  �Hn��N�  3�X�-@��mx�   npHy  ٬N�  3�X�".����fZHy  لN�  i|X�J�gHHy  مN�  h~X�-@���   �����f/N�  jX�/N�  jX�(J*L` ��p 0.������f�`� f�- e f� f�, f f� f�+ f f�$k ��    g� f�* f f�/N�  1�X�Hy  لHn��N�  ��P�Hy  ٬Hn��N�  ��P�/N�  1XX�Hy  لHn��N�  ��P�J�f �Z/N�  1�X�Hy  لN�  i|X�J�g �<Hy  مN�  h~X��   f �$Hy  ٬Hn��N�  ��P�J�f �/
N�  1�X�Hy  ٬Hn��N�  ��P�J�f ��Hn��N�  3�X�-@��m ���   n ��Hy  ٬N�  3�X�".����f ��Hy  لN�  i|X�J�g ��Hy  مN�  h~X�-@���   �f ��. _��g. 0��g. .��fN. L��fF/- /a tP�� | d Hy  ٬/a \P�� | f /N�  jX�/
N�  jX�` �/` �*y  �B`  f - e f  f  �, f f  � f  �+ f f  �/N�  1�X�Hy  لHn��N�  ��P�Hy  ٬Hn��N�  ��P�/N�  1XX�Hy  لHn��N�  ��P�J�f  �/N�  1�X�Hy  ٬Hn��N�  ��P�J�flHn��N�  3�X�-@��mZ�   nRHy  ٬N�  3�X�".����f<Hy  لN�  i|X�J�g*Hy  مN�  h~X�-@���  ������f/N�  jX�(K*L(m ��    g&l ��    f ��L�< `��N^NuNV��/*y  �B`  � f  �/N�  1�X�J�  �Xg0Hy  ��Hy  ٬N�  ��P�J�gHy  �Hy  ٬N�  ��P�J�fLHy  لN�  i|X�J�g:Hy  مN�  h~X�J�f(Hy  ٬N�  4.X������fHy  ٬/a NP�� *m ��    f �^*_N^NuNV��//J�  ��g �*y  �B` �- f f �/N�  1�X�Hy  لN�  i|X�J�g |Hy  مN�  h~X�-@���   m `Hy  �Hy  ٬N�  ��P�J�f F(m ��    g DH�H�_��   b  ��@0; N�  0� ��� � ������ � ����� � � �(l `�/N�  1�X�Hy  �Hy  ٬N�  ��P�J�fvY���Hy  لHy  �Hn��N�  �Z�� Hn��/a P�J���f/N�  jX�`2/.��Hy  �Hn��N�  �Z�� Hn��/a �P��   ��n� 
*l ` XHy  لa �X�J�fHy  ٬a �X�J�g �B*L` 0/N�  1XX�-|  ل�� .��R��� @ af� n�� 0m� R��� @ 7n� .��R��� @ @f� n��Jf�Y���9  مH�H�/ Hy  �Hn��N�  �Z�� Hn��/a  P�� | f J���g � /.��Hy  �$Hn��N�  �Z�� Hn��/a �P��   ��n �` �/N�  1�X�Hy  لa �X�J�f �Hy  ٬a �X�J�f �` �B/N�  1XX�Hy  لa lX�J�f ��` �" 
g �h g �`*m ��    f�(_*_N^NuNV��H�< `��*y  �B��    f �` - f f � 
f �, f f � f �+ f f �J� g �/N�  1�X�Hy  لN�  3�X�-@���   m ��   n �Hy  ٬N�  3�X�J�f t/N�  1�X�Hy  ٬N�  3�X�����f T/N�  1�X�Hy  لN�  3�X�J�f 6/.��Hy  �,Hn��N�  �Z�� Hn��/a hP�`  �- f f  
f , f f  � f  �J� g  �/N�  1�X�Hy  لN�  4.X�-@���   m  ��   n  �Hy  ٬N�  4.X�J�f  �/N�  1�X�Hy  ٬N�  4.X�����f  �/N�  1XX�9 a  لfp9 0  مff9 @  نf\J9  هfT/.��Hy  �5Hn��N�  �Z�� Hn��/a  �P�� B- /N�  jX�`$k ��    g* g � g ��*L(m ��    g&l ��    f�L�< `��N^NuNV��/*n Jg sf� pf�p`p *_N^NuNV��/*n J� g/- N�  ��X�/. N�  6X�+@ *_N^NuNV  a �a �a �a �N�  qNN�  rRaN^NuNV��H�8�`��*y  �B��    g �| `  �/a �X�`  ��    g�| `  �| `  �- f g
- e f  �/N�  1�X�Hy  ٬N�  4.X�. m  ��   n  �Hy  لa �X�J�gpHy  مa �X�J�f`//Hy  �|Hn��N�  �Z�� Hn��/N�  R�P�� | f *L(m ��    g �  g �L !g �R "g �J g �H f`- f fX/N�  1XX�Hy  لN�  3�X�. m<�   n4Hy  لHy  ƄHn��N�  �Z�� Hn��/N�  R�P�� &B- ` �lJ�  ܈g4 f./N�  1XX�9 _  لfHy  لN�  �DX�J�g� -` �0 f2/N�  1�X�Hy  لa �X�J�gHy  مa �X�J�f f �N f|  f f/a �X�/`  �&l ��    g  �J�  �Lgb f\ fV, d fN/N�  1XX�Hx Hy  ƊHy  لN�  ���� J�gHy  ƒHy  لN�  ��P�J�f/a jX�(M` �^ f �V f �NJf �HJ, f �@/a >X�/a 6X�L�8�`��N^NuNV��H�8�`��*y  �B��    f 	�` 	� f  �- f f  � f  �J, g,  g,  g
,  f  �J, f/N�  ��X�J�gl&m ��    g` f+ f g &fL/N�  1XX�Hy  لN�  3�X�. m0�   n(/N�  1�X�Hy  ٬N�  3�X���f/a TX�` 	$ f  � f  �- f f, f g$- e f, e g- d f  �, d f  �/N�  1�X�Hy  لN�  3�X�. m �Hy  ٬N�  3�X�, m �/N�  1�X�Hy  لN�  3�X�-@��m �Hy  ٬N�  3�X�-@��m x��f r����f j�   ��m
�   o V, e f�   ��l B/a fX�(M` 4 f � f �, f f �/N�  1�X�Hy  ٬N�  3�X�. m j�   n `Hy  لHn��N�  ��P�/N�  1�X�- f f  Hn��N�  4.X������f �Hy  لa PX�J�g �Hy  مa @X��   �f �Hy  ٬N�  3�X���f �Hy  ƜHn��a �P�J�g �� | f /Hy  ƟHn��N�  �Z�� Hn��/N�  R�P�� | d /Hn��Hy  ƣ` 0Hn��N�  4.X������f DHy  لa �X�J�g 2Hy  مa �X��   �f Hy  ٬N�  3�X���f Hy  ƪHn��a �P�J�g  �� | f /Hy  ƭHn��N�  �Z�� Hn��/N�  R�P�� | d /Hn��Hy  Ʊ`  �Hy  لa X�J�g  �Hy  مa �X��   �f  �Hy  ٬N�  3�X���fx� | f /Hy  ƸHn��N�  �Z�� Hn��/N�  R�P�� | d /Hn��Hy  ƼHn��N�  �Z�� Hn��/N�  R�P�` �- e g ��- d g �P- f f  �Hy  لa JX�J�g  �Hy  مa :X��  ��fnHy  ٬N�  3�X���f\Hy  ��Hn��a �P�J�gH� | f /Hy  ��Hn��N�  �Z�� Hn��/N�  R�P�� | e /Hn��Hy  ��` �0- e f  �Hy  لa �X�J�gnHy  مa �X��  ��fZHy  ٬N�  3�X���fH� | f /Hy  ��Hn��N�  �Z�� Hn��/N�  R�P�� | e /Hn��Hy  ��` �� f �- f f � f �, f f � f �+ f f �/N�  1�X�Hy  ٬N�  3�X�. m ��   n �Hy  لN�  3�X������f nHy  لHn��N�  ��P�/N�  1�X�Hy  ٬N�  3�X���f >Hy  لa �X�J�g ,Hy  مa xX��   f /N�  1�X�Hy  لa VX�J�g �Hy  مa FX��   �f �Hy  ٬N�  3�X���f �Hx Hn��N�  �2P�J�g �� | f /Hy  ��Hn��N�  �Z�� Hn��/N�  R�P�� | d /Hn��Hy  ��` P- e f p f h, f f ^ f V+ f f L/N�  1�X�Hy  ٬N�  3�X�. m .�   n $Hy  لN�  3�X������f Hy  لHn��N�  ��P�/N�  1�X�Hy  ٬N�  3�X���f  �Hy  لa X�J�g  �Hy  مa X��   f  �/N�  1�X�Hy  لa �X�J�g  �Hy  مa 
�X��   �f  �Hy  ٬N�  3�X���fn� | f /Hy  ��Hn��N�  �Z�� Hn��/N�  R�P�� | d /Hn��Hy  ��Hn��N�  �Z�� Hn��/N�  R�P�/` �� g �� f  �- f f  � f  �, f f  �/N�  1�X�Hy  ٬N�  3�X�. m  ��   n  �Hy  لHn��N�  ��P�/N�  1�X�Hy  لa 
�X�J�glHy  مa 	�X�-@���  ��nTJ�mPHy  ٬N�  3�X���f>Hy  ��Hn��a *P�J�g*| e /Hn��Hy  ��Hn��N�  �Z�� Hn��/` �� f  �- f f  � f  �, f f  �/N�  1�X�Hy  لa 
2X�J�g  �Hy  مa 	"X�-@���  �nlJ�mhHy  ٬N�  3�X�. mV�   nN/N�  1�X�Hy  لa 	�X�J�g4Hy  مa �X�-@���  �nJ�mHy  ٬N�  3�X���f| e *L(m ��    g&l ��    f �
L�8�`��N^NuNV��H�< `��*y  �B��    f �` � f $- e f  f , e f  g +f  �+  f  �J� g  �/N�  1�X�Hy  لa 	X�J�g "Hy  مa �X��   f Hy  ٬N�  3�X�-@���   m ��   n �/N�  1�X�Hy  لa �X�J�g �Hy  مa �X������f �Hy  ٬N�  3�X�����f �/a �X�/a �X�/+ /.��Hy  ��Hn��N�  �Z�� Hn��/N�  R�P�� ,| 
 (K f P- e f F f >, e f 4 f ,J+ f $J� g $k ��    g  f J* f  �J� g  �/N�  1�X�Hy  لa �X�J�g  �Hy  مa �X��   f  �Hy  ٬N�  3�X�-@���   m  ��   n  �/N�  1�X�Hy  لa fX�J�g  �Hy  مa VX������flHy  ٬N�  3�X�����fX/a �X�/a �X�/* /.��Hy  �Hn��N�  �Z�� Hn��/N�  R�P�� ,| 
 -k ��'j  %n�� (K*L(m ��    g&l ��    f �fL�< `��N^NuNV��//*y  �B��    g  � f  �- f f  �/N�  1�X�/a �X�. B���-n����B���`B .����  �< @-P��`(0�   gJ���g�J���fJ .����  �< @-P���R����   ��m�J���f*J���f$/a �X�`J���f/.��/a P�*m ` �FJ���f�/.��/.��/a *�� `�.*_N^NuNV��//B���-n����*y  �B��    g RH�H��   gHn�   gj�   g  ��   g  ��   g"�   g�   -g*m `�R���`�R���`�/N�  1�X�Hy  ٬Hy  لN�  ��P�J�f�/a �X�`�/N�  1�X�- f f�Hy  لa 
X�J�g�Hy  ٬N�  3�X��   m�Hy  مa �X�. ���� g ���� ���� f �d| e ` �Z- f f �P/N�  1�X�Hy  لa �X�J�g �4Hy  ٬N�  4.X�J�m � Hy  مa zX�. ���� g� ���� ���� g�` ��J�  �Xf,J���f  �J���f  �/9  �BHx Fa �P�. mt�   dll*y  �B`N/N�  1XX�Hx Hy  �>Hy  لN�  ���� J�gHy  �FHy  لN�  ��P�J�f$/a \X�`*m ��    g f�- d g�.*_N^NuNV��//*n a J�f$/. Hy  �PHn��N�  �Z�� /. Hy  �X`"/. Hy  �`Hn��N�  �Z�� /. Hy  �hHn��N�  �Z�� Hn��/N�  R�P�| f � N�  .$(@� | f B� B� Hn��/N�  R�P�B� 
)m   m !L +L )M (_*_N^NuNV��/*n aFJ�f/. Hy  �p`
/. Hy  �xHn��N�  �Z�� Hn��/N�  R�P�| f � *_N^NuNV  Hx Hy  ǀHy  ٬N�  ���� N^NuNV��H�8 `��*n (n &M/N�  3�X�J�l4`6�f�`, 0mB 7n< @f6 (f0S� )f(�f�| )��Bp`Jf�S� _g� .g� ag�p L�8 `��N^NuNV��/a �TJ�f&*|  ل #fV 0fP- x fH/a  �X�H�`HHx Hy  ǇHy  لN�  ���� J�gp�`&*|  ٬ #f 0f- x g�/. Hx SaP�*_N^NuNV��//*n `NJfF(m ��    g: .f4�. g
`* 9nR� 0l�  f =f  f
/aX�H�`*m ��    f�p�(_*_N^NuNV��//*n B���B��� -fR���R� 0f  �- x f  �T�`*�   alJ�   AmZ�   FnR .���Ї�   7-@��H�H�. �   0m��   9n� .���Ї�   0`��   fn� .���Ї�   W`�J�fJ���gH .��D�`Dp�`@H�H�. �   0m"�   9nr
 .��N�  �bЇ�   0-@��`�J�f�J���f� .��.*_N^NuNV��//*n  #fT -fR� 0fR- x fJT�H�H�. �   0m�   9o��   am�   fo��   Am�   Fo�J�gp ` 9nR� 0l�Jf�p.*_N^NuNV��//*n (m J� g/- N�  ��X�B�  m !L )m  +y  �( 
#�  �((_*_N^NuNuNV��H�<�`��*y  �B��    f �` � f �- f f |J� g t/N�  1�X�Hy  ٬N�  3�X�J�f V(m ��    g H f @, f f 6/N�  1�X�Hy  ٬N�  3�X�J�f &l ��    g 
 f + f f  �/N�  1�X�Hy  لN�  3�X�J�f  �Hy  ٬N�  4.X�J�f  �$k ��    g  � f  �J* g  �/
N�  1�X�9 a  لf9 0  مg  �Hy  ǐHy  ٬N�  ��P�J�fn/N�  1�X�Hy  لHy  ǔHn��N�  �Z�� Hn��/N�  R�P�/N�  1�X�Hy  لHy  ǚHn��N�  �Z�� Hn��/N�  R�P�/N�  jX�*m ��    f �h*y  �B`*L(m ��    f��  �Bg  f  �J- g  �/N�  1�X�Hy  لN�  3�X�J�fhHy  ٬N�  3�X�. �   mP�   nH(m ��    g< fJJ� gD&l `6 f, + �� f"$k ��    g"/
N�  ��X�J�f*m ` �\&k ��    f�(m ��  �Bg�H�H�_��   b��@0; N�  F��LL����������LLLL�������������������������� F(l `�/N�  1�X�Hy  ٬N�  3�X�, Hy  ٬N�  3�X�, �   m�   n��f�J�f �>9 #  لgf9 a  لg\9 _  لgR9 .  لf
9 L  مg>9 0  لm
9 9  لo*Hy  لN�  3�X�, �   m ���   n �Լ�g ��&m ��    fX`  �/N�  1�X�Hy  لN�  3�X�J�f  �Hy  ٬/Hy  ǠHn��N�  �Z�� Hn��/N�  R�P�&k ��    g^H�H��   g��   fH/N�  1�X�Hy  لN�  3�X�J�f  �Hy  ٬/Hy  ǧHn��N�  �Z�� Hn��/N�  R�P�(m ��  �Bg ��H�H�_��   b P�@0; N�  lD � �D � � � �DD � � � �DDDDDDDDDDDDD l(l `�Hy  ٬N�  3�X�J�f �~/Hy  لHy  Ǯ` �P/N�  1�X�Hy  ٬N�  3�X�J�f�/Hy  لHy  ǵHn��N�  �Z�� Hn��/N�  R�P�/N�  jX�*L` � /N�  1�X�Hy  ٬N�  3�X�J�f �b/Hy  لHy  ǼHn��N�  �Z�� Hn��/N�  R�P�` �4/N�  1XX�Hy  لN�  3�X�J�f �/Hy  ��Hn��N�  �Z�� `�H�H�/ Hy  ��Hy  μN�  �L�� ` �|/N�  1�X�9 _  لgH9 #  لg>9 .  لf
9 L  مg*Hy  لN�  3�X�, �   m �0�   n �&��g � Hy  ٬N�  3�X�, m ���f ��` �/N�  1�X�9 #  لgHy  لN�  3�X��   f ��Hy  ٬N�  3�X�, m ���   n ����f �,` ��/N�  1XX�Hy  لN�  3�X�, m ���   n ����f ��` �|L�<�`��N^NuNV��H�0�`��*y  �B��    f  �`  � f  � f  �, f f  �J, g  �/N�  1�X�Hy  ٬N�  4.X�J�f  �/N�  1�X�Hy  لN�  4.X�J�flHy  ٬N�  4.X�. �   mT�   nL/N�  1�X�/Hy  لHy  ��Hn��N�  �Z�� Hn��/N�  R�P�//N�  B�P�/N�  jX�(M*L(m ��    f �*L�0�`��N^NuNV��//J�  �Xf *y  �B��    f  �`  f  �- e f  � f  �, e f  �/N�  1�X�Hy  لHn��a  �P�Hy  ٬Hn��a  �P��   ��f  ��   ��f  �/N�  1�X�Hy  لHn��a  �P�Hy  ٬Hn��a  �P��   ��f\�   ��fR .������fH .�谮��f> .������f4 .�찮��f* .��T�����f .��T�����f| f /N�  jX�(M*L(m ��    f ��(_*_N^NuNV��H�0�`��*n (n *����� af: 0m4 7n. @f(Jf$*�    n ( H�H��   (+@ B� `  �(n  af  � 0m  � 7n  � @fz (ft~ -G�� -f*~R�`$ )g"r
 .��N�  �bH�H�Ё�   0-@��Jf� )f4Jf0*�    n ( H�H��   (+@ J�f .��` .��D�+@ L�0�`��N^NuNuNV��H�< `��*y  �B��    f 
�`  f �- f f � f �, f f � f �J+ g
+  f zJ+ f/a �X�J�g f/N�  1�X�9 a  لf
9 @  نg69 _  لg,9 .  لf
9 L  مg9 0  لm 9 9  لn Hy  ٬N�  3�X�J�f �/N�  1�X�Hy  ٬N�  3�X�J�f �Hy  لa 
@X�-@�������g �/N�  1�X�J���m �   ��nHx Hy  لa 
rP�J�f  ��   ��m�   ��nHx Hy  لa 
HP�J�fV�   ��m�   ��nHx Hy  لa 
 P�J�f.�   ��m :�   ��n .Hx  Hy  لa 	�P�J�g Hy  ل0.���   / Hy  ��Hn��N�  �Z�� Hn��/N�  R�P�� .B- /N�  jX�(K` 	 f �- e f � f �, f f � f �+ f f �$k ��    g � f �J* g
*  f zJ* f/
a �X�J�g f/N�  1�X�9 a  لf
9 @  نg69 _  لg,9 .  لf
9 L  مg9 0  لm 9 9  لn Hy  ٬N�  3�X�J�f  �/N�  1�X�Hy  ٬N�  3�X�J�f  �Hy  لa 6X�-@�������g  �/N�  1�X�J���m�   ��nHx Hy  لa hP�J�f,�   ��m  ��   ��n  �Hx  Hy  لa <P�J�gjHy  ل0.���   / Hy  ��Hn��N�  �Z�� Hn��/N�  R�P�� .B- /N�  jX�/N�  jX�(J` NJ�  �Xg �NJ�  �Xg �.J�  �Xf b f Z- e f P f H, f f > f 6J+ g
+  f &J+ f/a 
X�J�g /N�  1�X�9 a  لf
9 @  نg69 _  لg,9 .  لf
9 L  مg9 0  لm  �9 9  لn  �Hy  ٬N�  3�X�J�f  �/N�  1�X�Hy  ٬N�  3�X�J�f  �Hy  لa xX�-@�������gr/N�  1�X�J���m�   ��nHx Hy  لa �P�J�f(�   ��m:�   ��n0Hx  Hy  لa �P�J�gHy  ل0.���   / Hy  ��` �� f j- d f ` f X, e f N f F+ f f <$k ��    g . f &* f f -j ��g  n�� f J( g
(  f  � n��J( f/a `X�J�g  �/N�  1�X�9 a  لf
9 @  نg69 _  لg,9 .  لf
9 L  مg9 0  لm  �9 9  لn  �Hy  ٬N�  3�X�J�fv/
N�  1�X�Hy  ٬N�  3�X�J�fZHy  لa �X�-@�������gB/N�  1�X�J���m2�   ��n(Hx  Hy  لa P�J�gHy  ل/.��Hy  ��`  f &- d f  f , f f 
 f J+ g
+  f  �J+ f/a 4X�J�g  �/N�  1�X�9 a  لf
9 @  نg69 _  لg,9 .  لf
9 L  مg9 0  لm  �9 9  لn  �Hy  ٬N�  3�X�J�fv/N�  1�X�Hy  ٬N�  3�X�J�fZHy  لa �X�-@�������gB/N�  1�X�J���m2�   ��n(Hx  Hy  لa �P�J�gHy  ل/.��Hy  �` �� f  �- f f  � f  �, f f  � f  �J+ g
+  f  �J+ f/a X�J�g  �/N�  1�X�Hy  لN�  3�X�-@���   m^�   nVHy  ٬N�  3�X�J�fD/N�  1�X�Hy  ٬N�  3�X�J�f(Hy  لa �X�-@�������g/.��/ Hy  �` �" f  �- e f  � f  �, f f  � f  �+ f f  �$k ��    g  � f  �J* g
*  f  �J* f/
a X�J�g  �/N�  1�X�Hy  لN�  3�X�-@���   mf�   n^Hy  ٬N�  3�X�J�fL/N�  1�X�Hy  ٬N�  3�X�J�f0Hy  لa �X�-@�������g�   n/.��/ Hy  �` �� f `- d f V f N, e f D f <+ f f 2$k ��    g $ f * f f -j ��g  n�� f  �J( g
(  f  � n��J( f/a �X�J�g  �/N�  1�X�Hy  لN�  3�X�-@���   m  ��   n  �Hy  ٬N�  3�X�J�f  �/
N�  1�X�Hy  ٬N�  3�X�J�frHy  لa  �X�-@�������gZ�   nR/.��/ Hy  �Hn��N�  �Z�� Hn��/N�  R�P�� .B- /N�  jX�/N�  jX�/
N�  jX�(n��*L(m ��    g&l ��    f ��L�< `��N^NuNV��//. N�  i|X�J�gL-|   �� . R�/ N�  h~X�-@��~ ` .������g .���-@��R��    m� .������f `p�.N^NuNV��/*n  afL- @ fDV�Jf  ~J� g� ( . �   0�� )Bp`d )gR�Jf�JgRJ� g�� +`� _g .f- L g 0m, 9o`$R�Jf�J� g�� + . �   0�`� (g�p *_N^NuNV��//*n J- gp` �H�H�S��   %b ��@0; N� JJ�� �&� � ��� L L L L L� \ \ \ \ \�������&������ L*m ��    f�` H/N�  1�X�9 a  لf9 0  مg (9 a  ٬f�9 0  ٭f�` /N�  1�X�9 a  ٬f�9 0  ٭f�`  �/N�  1�X�Hy  لN�  4.X�J�g  �Hy  ٬N�  4.X�J�g ��9 a  لf9 0  مg  �9 a  ٬f �D9 0  ٭g  �` �4J- g  �` ��/N�  1XX�9 a  لf �9 0  مg\` �J� g ��(m ` f
 - �� g:(l ��    g ��J, g�` ��/N�  1XX�9 a  لf ��9 0  مf ��p (_*_N^NuNV��//*n J- gp` \H�H�S��   %b H�@0; N� ��<||<F �< � �<



 �< \ \ \ \ \<<<��<<�<<<<<<�*m ��    f�` �/N�  1�X�9 d  لf9 0  مg �9 d  ٬f�9 0  ٭f�` �/N�  1�X�9 d  ٬f�9 0  ٭f�` �/N�  1XX�9 d  لf�9 0  مf �xJ9  نf �n` ��/N�  1XX�9 d  لf �T9 0  مf �H` 4/N�  1�X�9 d  لf9 0  مg 9 d  ٬f �9 0  ٭f �`  �/N�  1�X�Hy  لN�  3�X�J�g  �Hy  ٬N�  3�X�J�f ��` �dJ- g  �` �X/N�  1�X�Hy  ٬N�  3�X�J�f ��` �6/N�  1XX�9 d  لf ��9 0  مgr` ��J� g �x(m `* f  - �� f(l ��    gD/a ��X�`<(l ��    g �>J, g�` �4/N�  1XX�9 d  لf �9 0  مf �p (_*_N^NuNV��H�8�`��*n A�� &HS�m - R�  @p `
/N�  ��X�. �   
g$�����fHx  Hx  /N�  ���� `  ��`�BA�� &H+ . f�Hx 	/Hy  �$N�  ���� J�f�Hk a  �X�. Hx Hx N�  �vP�(@��    f Hy  �.Hy  μN�  �LP�Hx��N�  �X�Hk N�  6X�(� ��  ܔ @)P  ��  ܔ @ �` �L�8�`��N^NuNV��//*n /a:X���  ܔ @(P`//N�  ��P�J�fp`(l ��    f�p (_*_N^NuNV��//*n ~ `H�H�V�"�.Jf�0�   ?.*_N^Nu /  o `  "L@  � Nu o  / `  L  �Nu /  o `  "L@  �Nu /  o `  "L@  � Nu o  / `  L   �Nu /  o `  "L@  �Nu / "/ `  LA Nu / "/ `  L Nu / "/ `  LA Nu / L/  Nu / "/ `  LA  Nu / "/ `  L  Nu / "/ `  LA  Nu / L/   NuNV��H� �`��*n ~ | `* 9nPr
 N�  �bH�H�Ё�   0. `.R�R�`(R�H�H��   	g��    g��   +g��   -g� 0l�J�g D�` L� �`��N^NuNV��H�8�`��*n ~ - �   @ f J� g - �� fJ�f- �   Df/N�  ��X�J�f8- H�H���  ϼ @&P(m  ��, n/N�  �X������f�p�`  �p `  �/Hx  /. /N�  ���� -@��g��S�, ��ݭ - H�H���  ϼ @ �� J�lr `"��l
/N�  �*X�ކJ���g$- �   Dg/N�  �X������g �v `ݮ ` �LL�8�`��N^NuNV��H�0�`��A�  . N�  �&/. N�  ��X�*@��    fp `(M . V�rN�  ��. `B�S�l� L�0�`��N^NuNV  /. N�  ��X�N^NuNV��H� �`��*n .. ,. -�� -   g  ��   lfJ� g`-  fX*(J�f$Hx Hx  - H�H�/ N�  �j�� "��؁`��- �   �fJ�o��n - �� ��m
٭ ��`  �-  g+m  -�� //- H�H�/ N�  �j�� ( B�`F- �   �g:/N�  ��X�-  gB�-�� +m  //- H�H�/ N�  �j�� ( �����fp�`p L� �`��N^NuNV��/A� -H��Hy  ή/.��/. N�  ���� . 9   κgp�` .N^NuNV��/A� -H��/. //. N�  ���� .  n (  gp�` .N^NuNV��H�0�`��*n (n .. ,. S�m�-��H�H���f� `p L�0�`��N^NuNV��H�8 `��*n A� &HJ� f
/N�  ��X�  f g  �  �   Dg*(|  Π`, �   @g
/N�  ��X��� ��  ϸe�+m   gp`- H�H���  ϼ @ �� / /- - H�H�/ N�  ���� *�S�m m p R� `$�����g   `  �   �g��B�p�L�8 `��N^NuNV��//*n (n ��g`Jfp `�g�H�H�S�H�H���(_*_N^NuNV  N�  �(/ /. /. a2�� N^NuNV��/*n /N�  �X�//. /. a
�� *_N^NuNV��H� �`��*n ��    gJ� g n Jfp `  � n ( + fp`p .  n H�H��   ag"�   rg,�   wf�J�gp`p �   `J�gp`p �  `
J�gp`p , Hx�//. N�  ���� * m �|B�E J�g <   �` n  rfp`p@ B� +m   L� �`��N^NuNV��/*|  Π`��  ϸep `�� - �   �f� *_N^NuNV��//A���*H*����+n  +m  |  |  A� -H��///. N�  ���� .  m B .*_N^NuNV�H�<�`�*n (n B���B.�[&M`
�   %gR�H�H�. f� ��-@�2gtѮ���   f,S�mp ", R�  A�p `N/p / N�  ��P�`<,  f/.�2//, N�  ���� Ю�2)@ `//.�2Hx /N�  ���� J�f,  gp�` F .��` >B���-n����-n����-n����-n����`f�   *f|X�  n -h����J���l .��D�-@��R���R� .g "J���g  � .��`  �R���`�   #g,�   +g��   -f�R���R�H�H�. �    f�R���`�R���`��   0fR���B���H�H�. �  ̹ @�   g �~r
 .��N�  �b"�   0Ё-@��R�`�p�-@��B���H�H��   hg  ��   lg  �-|  ˄�`A��[-H�\B���-n����H�H�. �   cg (n ��   Fg Nn j�    g ���   Dgv�   Eg G�e` R� *fX�  n -h����R�` �fB���H�H�. �  ̹ @�   g �Fr
 .��N�  �b"�   0Ё-@��R�`�R���R�` �<~d-|   �.R���` -|   �.`R���-|   �.`-|   �.J���l-|   ��J���g `(-|  ˅�`��   �RgP .�RD�-@�R`D�   df  X�  n -h���R�   df$J��Rm�J���g
-|  ˇ�``J���g-|  ˉ�`�   Xf <  ˋ` <  ˜-@�:A��p&H$K`F0.�T�   -@�* .�R�����-@�R".�.N�  �t�Ю�:Ю�* @S��A��R .�.N�  ��J��Rf� ��Ю��-@��J���g��g �   Xgb�   og<�   xgHJ���lB���J���lB��� 
��-@�2Ю��Ю�� n�`Jf �r ` ��   ��l�-|   ��`�-|  ˭�``�-|  ˰�``�J���l-|   ��J���gP�  n -h���J-h���F`X�  n -h���NJ���g6Hn�>Hn�B .��R��   l .��R�`p/ /.�J/.�FN�  ���� `0Hn�>Hn�B .��R��   l .��R�`p/ /.�NN�  ���� &@J��>g
-|  ˳�``J���g
-|  ˵�``J���g-|  ˷�`A��e$HJgH�H�`p0�J���fJ���g� .-n����`
Jg�S���J���n�A��e&HJ���g
".�J .�F`
 .�NN�  �&/9  �p/9  �l// N�  ���� gR .�BS�-@�2J�l0D�-@�2`(r
 .�2N�  �t�   0S��\ n�\�A��2p
N�  ��J��2g`�S��\ n�\� 0A��Y .�\��b�J��Bn6J���g
".�J .�F`
 .�NN�  �&/9  �x/9  �t// N�  ���� fp+`p-S��\ n�\� �  ̹ @  gpE`peS��\ n�\�` ��J���l-|   ��J���gP�  n -h���J-h���F`X�  n -h���NJ���g0Hn�>Hn�B�   <��l .��`p</ /.�J/.�FN�  ���� `*Hn�>Hn�B�   <��l .��`p</ /.�NN�  ���� &@J��>g .��D�".�B��o 0g
-|  ˹�``J���g
-|  ˻�``J���g-|  ˽�`A��e$H-n�B�2B��6J��2oJg
�   �6mp0`
R��6H�H��S��2n�J���fJ���o� .�   <��l .��`p<-@�2 .�����2-@��`$R��BoJg
�   �6mp0`
R��6H�H��S��2l�A��e&H` �J���l-|   ��J���gP�  n -h���J-h���F`X�  n -h���NJ���g0Hn�>Hn�B�   ��l .��`p/ /.�J/.�FN�  ���� `*Hn�>Hn�B�   ��l .��`p/ /.�NN�  ���� &@J���g
".�J .�F`
 .�NN�  �&/9  ˀ/9  �|// N�  ���� f-|   �B-n���6J���f8/N�  ��X�-@�2���6l-@�6` .�6S�Ћ @ 0fS��6�   �6l�������Bm
 .�B����o .�6S�-@��` �� .�6���B-@��` ��X�  n  (��@�eA��e&HA� $H` ��X�  n &h��$KJ���l/N�  ��X���` �zJgS���l�S�` �j�   Gg �V�   Og �(�   Ug ��   Xg �"` ���   gg �*n"�   dg ���   eg �z�   fg ��` �\�   og ���   sg �`�   ug ���   xg ��` �0 n�`J( fr`rЁA��[���\Ј-@�6 .�����6n .�6Ѯ��J���g(`t , R�  @�  p `S�l�/Hx  N�  ��P�S��� .�����6l�`> .�`R��` @p ", R�  A�p `S�l�/ .�`R��` @p / N�  ��P� n�`Jf�`& , R�  @� 0p `S�l�/Hx 0N�  ��P�S���l�J��2o  ��   �2f$S�mp ", R�  A�p `j/p / `X,  f/.�2//, N�  ���� Ю�2)@ `://.�2Hx /N�  ���� `" , R�  @� 0`�S�l�/Hx 0N�  ��P�S���l�`> .�\R��\ @p ", R�  A�p `S�l�/ .�\R��\ @p / N�  ��P� n�\Jg`� , R�  @�  p S��� .�����6m �*S�l�/Hx  N�  ��P�`�L�<�`�N^NuNV  Hx  /. /. /. /. /. a.�� N^NuNV  Hx /. /. /. /. /. a�� N^NuNV��H�<�`��*n (|  �� . Ќ&@0. �  ��@�f2 . � ��J�fJ� gHx`Hx Hx 	N�  �<P�-A -@ /9  �/9  �/. /. N�  ���� lp`p  n  �g".  . @ -A -@ B9  ��B�/9  �/9  �/. /. N�  ���� g $|  � R�/9  �l/9  �h/. /. N�  ���� l  �/9  �t/9  �p/. /. N�  ���� m :-y  �|��-y  �x��/.��/.��/9  ̄/9  ̀N�  ���� -A��-@��/. /. // N�  ���� nR-n����-n����`�A� "*  N�  �� * ѕ/* //. /. N�  ���� l� J�� �    n�` /.��/.��/. /. N�  ���� N�  �@. �   0�A� -H��/.��/.�� N�  �// N�  ����  n��N�  ��R�/9  ̌/9  ̈/.��/.��N�  ���� o  �A���"9  ̔ 9  ̐N�  ��` �j/9  ̜/9  ̘/. /. N�  ���� l\/* //. /. N�  ���� /9  ̤/9  ̠// N�  ���� lA� "*  N�  �� * ��`� J�� �    n�J� g�շ�  ��e  Է�  �c&|  �/9  ̬/9  ̨/. /. N�  ���� g��  ��e� 0`X".  . N�  �@. �   0� N�  �// /. /. N�  ���� // /9  ̴/9  ̰N�  ���� -A -@ ��e$(K 5m0��  ��f� 1  ��R�J� gR�`R�` �N� 0S�R 9n�B <  ��L�<�`��N^NuNV  Hx  /. /. /. /. a*�� N^NuNV  Hx /. /. /. /. a�� N^NuNV��H�<�`��*n (|  ͼ . Ќ&@0. �  ��@ �f( . � ��J�gHx`Hx Hx 	N�  ��P�-@ "9  � . N�  �lp`p  n  �g . @ -@ B9  ͼB�"9  � . N�  �g 8$|  �R�"9  �D . N�  �l."9  �H . N�  �m  �.9  �L`4A�  N�  �X * ѕ" . N�  �l� JP��    n�`  �." 9  �PN�  �l, ". N�  �o�" . N�  ��N�  ��* �   0�A� -H�� N�  ��"N�  �l n��N�  �:R�"9  �T N�  �o`"9  �X N�  ��. `�"9  �\ . N�  �m`:A�  N�  �J * ��" . N�  �l"9  �`N�  �m� JP��    n�J� g�շ�  ͼe  ʷ�  �
c&|  �
"9  �d . N�  �g��  ��e� 0`\ . N�  ��. �   0� N�  �//  . N�  �&// N�  ���� // /9  �l/9  �hN�  ���� N�  �R-@ ��e$(K 5m0��  ͼf� 1  ͼR�J� gR�`R�` �X� 0S�R 9n�B <  ͼL�<�`��N^Nu"/  / @ NuL�  `L�  A 3�   �p`3�   �pH�> �U��Uð�c�A�C��B�BD fJ�g  zJf�fҀ�`l��`h< �< � �gl<�DF mQF��f�쨴fҀd&�REE �m`  ���kgt�[���SEngBE���   �d
�REE �gT����� L� |3�   �pNu�J�g <  `�fִg� <  "`  / ?9  �pBgN�  ��P�" `�B�`� <   `�L�    g��   fB�`��� e
`B�� l: g��   fB�`��� d  g�A`�� l��< NuB�" `/<   //<  /<   N�  ��P�"J�f��A`�o  3�   �r`3�   �rH�? L�  �U��UŰ�c�B�C�EH��a JGf( ��gx��JFf
��`0� F�gj� �FDGQGm ����f�J�f�`^Gk��Q���JkցՀd��RFF�m`^����dFED�@�a �a �M� "L� �Nu� a `�(��g <  `�FJj� <  "`  / ?9  �rBgN�  �<P�`� <   `�H�� L�  (Ȁk ��   fJ�fB�`��   fJ�fB�`�B�C��f(��g�< 
< L� NuL�  H�< �� ���BCBD @� A� RSDoBR RSCofR�蘘C6HA��4 ��B@��䀁�H�H�HB�Ђ�D a H����L� <Nuf
SD�b�RD`��fJ�fJ�f"<  B`ZJ�g2"<  `NgJ�f�B�`�J�g
SC�d�RC`�"<   J�f,"<  A`$ <   �`���eJ�g�@���`p ��  ` ��//<   N�  ��P�` �nH�? L�  * ���グ�c�B�Ca �:,�GE�g  �JGg  �� � H�� L� :/ ��������B�:/ �� 
օӇ:/ �� օӇ:�� օӇ:/ �� 
ԅч:�� ԅчH@:�� 
҅�GH@�� 6HCBAHAւчЁ$ F�a ��� "L� �Nu�  �g"<   `$*�G����g"<  `J�f J�f"<  0`  / ?< BgN�  �<P�`�<<�a �`�. ��gSF��j�RF` �$<� `�B�B�` �� / " H�> a �` / H�> " a �a  �L� |NuL�  H�8 aa �`L�  H�8 aa � L� Nu$<��  & HCĀ��(���f< J�g,< `&HB�JB�f4<` < J�g< `� SB< B2Nu m��� ���  `B>�B�F�Ca>ap,  �A�K�Nux����,<  �.̂��(ȃ��⊄�(΀��ȁ��∀�NuJ�fF  mF  �BJ�gk��[���Z� Nu<<�RNuJ�kSF��JFnF��mJDF��Q���BF�   d
R�d��RFF�l,(<��� ƄȂ����$�eF�gBFx軄F�NuB�B�Nu$<��  B�NuH�? L�  L�  $3�   �t* ��B�a^:�G8< a L,8< a BᏄ�g� ��$&<F�a �B` �. � ��HG�O�DfJ�fJ�gRGSG��  g�Nu8<��@�Aa��B�C�Fg�Dg� a�g&�Dg  �� ��Nua�J�k2�FgJJ�g "<  `PJ�k2��f"<  A`@"<   `8$<��  `  �J�f"<  R`""<  `"<  Q`J�f�J�f�"<  B`  X�/?9  �tBgN�  �<P�`  �J�g"<  `�J�j4XO`  ��Gf��l<$ HB�N�FHB����  b$<�� J�jT�B�`B�B�XO`dB�փՂ��\���	ǖ���[���jցՀ	�JD]���NuH�? L�  L�  $3�   �t*x�a ��8SG�Go
��<SFa�F a ��a ���� "L� �Nu"/ H�   �va`   o HB4H� L�   �vNu&HC��BBf< J�g*< `$ �f4<` B< J�g< `< SB< B ����B�Nu o L� 6HB o NuH�   �va�a �L�   �vNu8 m�� ��  �`*J�g
 PD����f� gkSD�j�D �a(  �g
��" �K�Nu/<   /<   N�  ��P�" NuJ�kSD�JDnD��m"DR�BD�   �d�RDD �l�U��NuB�Nu <   �Nu / H�8 " a$a �V L� Nu / H�8 " a ��a L� NuBBvJ�jD�� B�Nu la*�BJ�fJ�kJCjD�Nu/<  p/<   N�  ��P�" Nux JBk&�Dm
J�fD�D�@`���x�S�$ Ąf.ȁ����`$DB�Dm" B��D`�x�S�F�Ȁ������ B�NuH�^ "/  / �U����BCBD RSCo^< RSDoZ< �䙖Dm0Ѐ��[���Z� `ЀЁZ���[���jЁ�kg�[���Z� `�C�a ������/@ L� zNuf*�`�fSD�b�f"<  Q`(RD`��   �g�"<  `"<  �   �f"<  R//<   N�  ��P�`�L�  H�< * ���ば�c�A��BD BC�C �g>J gz< �< �4 6H@HA������ւ�C HCЃD ~a ������L� <Nu �g"<   `BJ�g"<  `
J�f"<  0//<   N�  ��P�`�< � `�J�g�k�SD�j�` �~ <� `�B�`�"/a �� _ �Nu"/�Aa � _ �Nu"/a � _ �Nu"/�Aa �� _ �Nu/Hy  �|H�? $&` �: _ � �Nu/Hy  ��H�? $ &B  "` � _ � �Nu/Hy  ��H�? $&` �. _ � �Nu/Hy  ��H�? $&` �� _ � �NuNV  3�   ݢ�   ݠ�    fp `p�  ݡ�   
 g
#�  Έ  ݘHx N�  ��/ N�  �xP� 9  ݘN^NuNV  3�   ݢ�   ݠ�   ݡ�   
 g#�  ΐ  ݜ#�  Ό  ݘHx N�  ��/ N�  �xP�"9  ݜ 9  ݘN^NuNV��H�8�`��.. ,. *n J�o  �J�o  �- �   @ f J� g - �� fJ�f- �   Df/N�  ��X�J�fV- H�H���  ϼ @&P" N�  �b* (m  ��( n./N�  �X������f� ЇS�"N�  ��"�� `  �p `z��d ` ( //. /N�  ���� ��٭ - H�H���  ϼ @ �� J�lr `"��l
/N�  �*X���f- �   Dg
/N�  �X� `ٮ ` �NL�8�`��N^NuNV��/*|  Π`
/aX��� ��  ϸe�*_N^NuNV��//*n ~���    gj- �   �g:- �   gp `/aTX�. - H�H�/ N�  �X�J�l~�#�     h-  g/- N�  ��X�B� B- B�+m   .*_N^NuNV��/*n - �   fB�`6-  f"-  gJ� g - �� c
/a RX�`�-  gp�`p *_N^NuNV��/*n - �   R@ Bf|- H�H���  ϼ @ - ��d  �R�  @�   
f  �/a  �X������g6`  �n ��Hx Hn��- H�H�/ N�  �"�� �   g  � -   p�`  �- �   @ g�- �   @ f J� g - �� fJ�f- �   Df/a X�J�f�- �   Df �/aDX�S�mp . "- R�  A�p `/p . / a ��P�-  f �fp . *_N^NuNV��H�0�`��*n (m  - ��. +L - �   Dgp `- H�H���  ϼ @ �� *�- H�H���  ϼ @ �� J�lr `"��l/a �X�J�o( / /- H�H�/ N�  �"�� ��g
 -   p�`p L�0�`��N^NuNV��/*n - �   @ g*- �   �fp�`  �- H�H������ �   @ J� f/ahX� - �� fT- �   DfH- H�H���  ϼ @ �� *�- H�H���  ϼ @ �� J�lr `"��l/a  �X�p *_N^NuNV��//*n - H�H�. �   l$ ��  Θ @+P ` -   - �   `&HxN�  ��X�+@ f� ��  ݤ+@ �    - H�H���  ϼ A �+m  /N�  �(X�J�g-  f - @ .*_N^NuNV��//*n - H�H���  ϼ @ �� . l- H�H���  ϼ @+P `��l*�.*_N^Nup% o "/ N@ep NuN�  �<NV��H�8�`��*n (n .. &M`�S�l� L�8�`��N^NupN@NuNV��//*n A� (HJf� ��(_*_N^NuNV��H�8�`��J�  �f8 <  � �   #�  � <  � �   #�  �#�  �  \#�  �  X . ^���. *y  X 9  ��"9  �����nx �����&@-   fX(U,   fD*�X�  �S�  ���f�(U "҇��m> Ї#�  X��c  � @#�  ` @ �Y�  �`  � "҇��l� �����*@��f� � �� �  @ `$J�  Tfp `  � y  TN�0�  � �   #�  � / N�  ��X�(@ �����g� y  \ � 9  \X���g y  \  �    � й  � Y�(�#�  \ <  � �    y  \ � 9  � Q�ѹ  �T�  �` ��S�  � 9  X �   *� Y���  �A�  L�8�`��N^NuNV��//*n (MY�#�  X �����(�"��Y�ѹ  �R�  �(_*_N^NuNV��H�<�`��*n -  ��g/a�X� -��"���. /. a ��X�(@��    gJ��gF&M$L . V��, ��d.`$� S�J�f���d" �Ќ��e "�Ё"��"Ҁ A �  ` L�<�`��N^Nu 9  �$ѯ p o N@e 9  �$#�   �$NuN�  �<p o N@e�#�   �$p NuNV��H�0�`��*n (n .. ��g`�fJfp `S�l�J�m�H�H�S�H�H���L�0�`��N^Nup o N@ep NuN�  �<NV��Hn��HxT/. N�  �P�� J�lp `pN^Nup6 o "/ "o N@eNuN�  �<p o "/ "o N@eNuN�  �<p o "/ "o N@eNuN�  �<p o "/ "o N@eNuN�  �<NV��H�8 `��*n (n &MJf�S��f� L�8 `��N^NuNV��H�8 `��*n (n &M�f� L�8 `��N^Nup
 o N@ep NuN�  �<p o "/ "o N@eNuN�  �<#�  hp�NuNV  N�  ��/. N�  �`X�N^Nup o N@Nr  (C) Copyright 1983 UniSoft Corp. Version III.1.4  UniSoft Systems usage:c2 [-KPSdls] [if [of] ]
 r c2: can't find %s
 w c2: can't create %s
 iterate
 comjump
 rmove
 | end output: t->op=%d, t->subop=%d, t->code=%d, t->labno=%d, t->misc=%d
 .L%d: 	| line %d 	| line %d output: opcode = %d
 	.L%d%s 	| line %d 	| line %d 	.L%d 	| line %d 	| line %d c2:out of string storage space
 %d iterations
 %d jumps to jumps
 %d inst. after jumps
 %d jumps to .+2
 %d redundant labels
 %d cross-jumps
 %d code motions
 %d branches reversed
 %d redundant moves
 %d simplified addresses
 %d loops inverted
 %d redundant jumps
 %d common seqs before jmp's
 %d skips over jumps
 %d redundant tst's
    	  N                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 ��0x1044 %d: %s  -
 #0 #0 c2:out of node storage space
                                                                                   #0  %s,a0 %s,a0 %s,a%d %s,a%d %s,a%d %s,a%d sp@- %s,a0 a0@ sp@- %s,a0 a0@ a%d,%s c2: Ax byte optimization error on '%s'
 #%d,%s #0x%lx,%s a%d,d0 a%d,d0 sp@- sp@ sp sp@- %s,sp@ #%ld,sp a%c,sp@ #%ld,sp d%d,sp@- a%d@     �  �  �  �  �  �  �   �#  �&  �)  �,  �/  �2  �5  �8  �;a%d,a%d #0,%s sp@(-.M sp@(-132) +3 d%d %s,d%d +1 d%d %s,d%d d%d %s,d%d +2 d%d %s,d%d d%d %s,d%d d%d %s,d%d d%d %s,d%d +2 %s,d%d d%d,.L%d d%d,.L%d d0 d1 d2 d3 d4 d5 d6 d7 a0 a1 a2 a3 a4 a5 a6 a7 sp@(-.M sp@(-132) %s,sp@- %s,sp@- sp@+,%s sp@+,%s %s,sp@- sp@+,%s a6@(-. a6@(-.   a0@ %s,a0 %s,a0 d%d,%s d%d,%s %s,d%d %s,d%d %s,d%d d%d c2:dregopt error: op=%d
 %s,a%d  #%d,%s #%d,%s #%d,%s #%d,%s #%d,%s #%d,d%d #%d,d%d #%d,d%d  	.globl	_ c2:out of global name storage space
    �T     �X     �\    �`    �d    �h    �l    �p    �t    �x    �|  	  ʀ  
+  ʄ   +  ʈ  +  ʌ  +  ʐ  +  ʔ  +  ʘ  +  ʜ  +  ʠ  +  ʤ  +  ʨ  	+  ʬ  
,  ʱ     ʵ     ʼ   %  ��     ��     ��   	  ��   
  ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     �      �     �     �   '  �   (  �   )  �   *  �     �$     �(   -  �,     �0     �4   .  �9     �?   &  �E     �J     �O      �U   !  �[   "  �`   #  �f   $        bra beq bne ble bge blt bgt bcs bhi bls bcc jra jeq jne jle jge jlt jgt jcs jhi jls jcc dbra jmp .globl .word mov clr not addq subq neg tst asr asl lsr lsl ext cmp add sub and or eor muls mulu divs divu jbsr jsr bsr lea pea btst movem moveq link unlk .text .data .bss .even .end                           - +   0123456789ABCDEF 0123456789abcdef 0x 0X - +   - +                                                                                                    F����n    CA�y7��    A�ׄ       @È        @Y         @$         C@      @$      @$      @$      @$      @$      ?�      @$              @$                (((((                  H����������������������                                                                                                                                                                                                                            t�Ů    Z�   L��    F@    B�     A      K�  A   A   A   A   A   ?�  A       @$                                              �L  �D                               ��  ��                                                                                                                                                                                                                                                ϸ          �                                                                                              l